
/*************************************************************************/
// Full Adder Structural Code using cells from OpenRoad's nangate45 lib 
/*************************************************************************/

# clock Path - Clock - > CLK ...mlb .

module fulladder (A,B,C,Sum,Carry,Clock, Scan_clk,Scan_en,cg_en, gen_clk_mux );

input A,B,C,Clock,Scan_clk,Scan_en,cg_en, gen_clk_mux;
output Sum,Carry;
wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;
endmodule

module fulladder (B,C,a,SUM,A, Carry,Scan_clk);
input A,B,C;
output SUM,Carry,Scan_clk;
wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;
endmodule


module fulladder2 
input a,inpu, b;
output x,z;
wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;

endmodule

module fulladder3
input a ,b;
output x,z;
wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;
endmodule

module fulladder4 
input a ,65;
output x,z;

//Full Adder Structural Code using cells from OpenRoad's nangate45 lib

wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;
endmodule

