module fulladder (A,B,C,Sum,Carry,Clock, Scan_clk,Scan_en,cg_en, gen_clk_mux );
input A,B,C,Clock,Scan_clk,Scan_en,cg_en, gen_clk_mux;
output Sum,Carry;
wire  n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, CLK, mux_clock,gated_clock;
endmodule
